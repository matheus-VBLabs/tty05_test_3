

//IMPORTED BLOCK:AND2b
module AND2b( 
A, 
B, 
Y 
); 

//-----------Input Ports--------------- 
input A,B; 

//-----------Output Ports--------------- 
output Y; 

//-------------Code Start----------------- 
assign Y = A & B; 

endmodule




//IMPORTED BLOCK:inverterC
module inverterC( 
A,
Q
); 

//-----------Input Ports--------------- 
input A;

//-----------Output Ports--------------- 
output Q; 

//-------------Code Start----------------- 
assign Q = ! A;

endmodule




//IMPORTED BLOCK:one_hz_clock
`define clock_frequnecy 27_000_000
module one_hz_clock #(parameter DELAY = 1000)(input clk,            // clk input
								output reg out);  // output pin

  localparam TICKS = DELAY * (`clock_frequnecy / 2000);

  reg [26:0] counter = 0;
  
  initial out = 1;
  
    always @(posedge clk) begin
    	counter <= counter + 1'b1;
    	if (counter == TICKS) begin
    		out <= ~out;
    		counter <= 27'b0;
    	end
    end
endmodule




//IMPORTED BLOCK:counter_6bits
module counter_6bits(input in, output reg a, output reg b, output reg c, output reg d, output reg e,output reg f);
  reg [5:0] count;
  always @(posedge in)begin
    count <= count + 1;
    a <= count[0];
    b <= count[1];
    c <= count[2];
    d <= count[3];
    e <= count[4];
    f <= count[5];
  end
endmodule



//IMPORTED BLOCK:tune
module tune
(
    input clk, 
    input [9:0] freq,
    output reg out
)

;
    reg [20:0] aux = (13513513/freq);
    reg [20:0] count_freq = 0;
 
    
    initial begin
        count_freq = 0;
    end 

    always @(posedge clk) begin
        count_freq <= count_freq + 1;
        out <= 1;
        if(count_freq >= aux) begin
            out <= 0;
            if( count_freq == aux*2)
                count_freq <=0;
        end
    end


endmodule



// Automatically generated by ChipInventor Cloud EDA Tool - 2.1
// Careful: this file (hdl.v) will be automatically replaced when you ask
// to generate code from BLOCKS buttons.
module tt_um_chip_inventor_music__6_bit_count (
    input  wire [7:0] ui_in,    // Dedicated inputs - connected to the input switches
    output wire [7:0] uo_out,   // Dedicated outputs - connected to the 7 segment display
    input  wire [7:0] uio_in,   // IOs: Bidirectional Input path
    output wire [7:0] uio_out,  // IOs: Bidirectional Output path
    output wire [7:0] uio_oe,   // IOs: Bidirectional Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  wire btn1;
  wire buzzer;
  wire l1;
  wire l2;
  wire l3;
  wire l4;
  wire led0;
  wire led1;

 assign btn1 = ui_in[0];


 assign uo_out[0] = buzzer;

 assign uo_out[1] = l1;
 assign uo_out[2] = l2;
 assign uo_out[3] = l3;
 assign uo_out[4] = l4;
 assign uo_out[5] = led0;
 assign uo_out[6] = led1;

 assign uio_oe = 8'b11111111;

 assign uio_out = 8'b0;

 assign uo_out[7] = 1'b0;



//Internal Wires
 wire w_1;
 wire w_2;
 wire w_3;
 wire w_4;
 wire w_5;
 wire w_6;
 wire w_7;
 wire w_8;

//Instances os Modules
tune blk202_1 (
         .clk (clk),
         .freq (10'd264),
         .out (w_1)
     );

AND2b blk2_4 (
         .B (btn1),
         .Y (buzzer),
         .A (w_1)
     );

counter_6bits blk173_7 (
         .in (w_2),
         .a (w_3),
         .b (w_4),
         .c (w_5),
         .d (w_6),
         .e (w_7),
         .f (w_8)
     );

one_hz_clock blk80_8 (
         .clk (clk),
         .out (w_2)
     );

inverterC blk5_9 (
         .Q (l1),
         .A (w_3)
     );

inverterC blk5_10 (
         .Q (l2),
         .A (w_4)
     );

inverterC blk5_11 (
         .Q (l3),
         .A (w_5)
     );

inverterC blk5_12 (
         .Q (l4),
         .A (w_6)
     );

inverterC blk5_13 (
         .Q (led0),
         .A (w_7)
     );

inverterC blk5_14 (
         .Q (led1),
         .A (w_8)
     );


endmodule
