

//IMPORTED BLOCK:AND2b
module AND2b( 
A, 
B, 
Y 
); 

//-----------Input Ports--------------- 
input A,B; 

//-----------Output Ports--------------- 
output Y; 

//-------------Code Start----------------- 
assign Y = A & B; 

endmodule




//IMPORTED BLOCK:OR2b
module OR2b (a, b, y);

//-----------Input Ports---------------- 
    input a,b; 

//-----------Output Ports--------------- 
    output y; 

//-------------Code Start--------------- 
    assign y = a | b;

endmodule



//IMPORTED BLOCK:tune
module tune
(
    input clk, 
    input [9:0] freq,
    output reg out
)

;
    reg [20:0] aux = (13513513/freq);
    reg [20:0] count_freq = 0;
 
    
    initial begin
        count_freq = 0;
    end 

    always @(posedge clk) begin
        count_freq <= count_freq + 1;
        out <= 1;
        if(count_freq >= aux) begin
            out <= 0;
            if( count_freq == aux*2)
                count_freq <=0;
        end
    end


endmodule



// Automatically generated by ChipInventor Cloud EDA Tool - 2.1
// Careful: this file (hdl.v) will be automatically replaced when you ask
// to generate code from BLOCKS buttons.
module tt_um_chip_inventor_music__6_bit_count (
    input  wire [7:0] ui_in,    // Dedicated inputs - connected to the input switches
    output wire [7:0] uo_out,   // Dedicated outputs - connected to the 7 segment display
    input  wire [7:0] uio_in,   // IOs: Bidirectional Input path
    output wire [7:0] uio_out,  // IOs: Bidirectional Output path
    output wire [7:0] uio_oe,   // IOs: Bidirectional Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  wire clk;
  wire buzzer;
  wire btn1;
  wire btn2;
  
assign btn1 = ui_in[0];
 assign btn2 = ui_in[1];

 assign uo_out[0] = buzzer;

 assign uio_oe = 8'b11111111;

 assign uio_out = 8'b0;

 assign uo_out[7:1] = 7'b0;

//Internal Wires
 wire w_1;
 wire w_2;
 wire w_3;
 wire w_4;

//Instances os Modules
tune blk202_1 (
         .clk (clk),
         .freq (10'd264),
         .out (w_1)
     );

AND2b blk2_4 (
         .B (btn1),
         .A (w_1),
         .Y (w_2)
     );

tune blk202_7 (
         .clk (clk),
         .freq (10'd300),
         .out (w_3)
     );

AND2b blk2_9 (
         .B (btn2),
         .A (w_3),
         .Y (w_4)
     );

OR2b blk10_11 (
         .y (buzzer),
         .a (w_2),
         .b (w_4)
     );


endmodule
